module multiply(i1,i2,out4);
   input [15:0] i1,i2;
   output [31:0] out4;

   assign out4 = i1*i2;

endmodule
